`include "RBLWE.v"
`timescale 1ns / 1ps

module Testbench;

	parameter CLOCK_PERIOD = 10;
	parameter ITERATION_SIZE = 5;

	// Inputs
	reg clk,reset;
	reg load;
	reg start;
	reg [7:0]c1_in;
	reg [7:0]c2_in;
	reg r2_in;

	// Outputs
	wire message_out;
	wire valid;
	
	// Instantiate the Unit Under Test (UUT)

	RBLWE dut (
		.clk(clk),     //clock signal
		.reset(reset), //global reset signal
		.load(load),   //load input signal
		.c1_in(c1_in), //c1 coefficient input (one coefficient at a time)
		.c2_in(c2_in), //c2 coefficient input (one coefficient at a time)
		.r2_in(r2_in), //r2 coefficient input (one coefficient at a time)
        .start(start), //start signal (active one cycle)
		.message_out(message_out), //message output (one bit at a time)
		.valid(valid) //output ready signal (high if an output is available)
	);
	
	
	reg [2047:0] c1 [ITERATION_SIZE-1:0];						  
	reg [2047:0] c2 [ITERATION_SIZE-1:0];									 
	reg [255:0] r2 [ITERATION_SIZE-1:0];
	reg [255:0] m [ITERATION_SIZE-1:0];

	
	reg [2047:0] c1_temp;						  
	reg [2047:0] c2_temp;									 
	reg [255:0] r2_temp;
	
	integer i;
	integer j;
	
	initial begin
		//TEST VECTOR INPUT 0
		c1[0] = 2048'hABD2CD28588EDE0CD8C7E3686229C1253764BF347B1DAA1EC369F2671D3AE1FA08929B4F4B785D6AA8F5F7CF6536989719F258CE16A9129A1C03FF4DC368D50645E9DECBB75CA8057CF7DB12E21C28BD4EEE18D22A2AD124C3BB8D80C4CCCD65AB3D005DEB7FC949BEA0F0823D9E1CED76117DC2549E028589199DDC07AEAB53A2B53416389C36A42ACE51B277E288D07FABE78D45A344EF21E5D5349957C109512DD9A7C1B5F0D757A9844D0834E7CBDCCD7EC02E018E04396E809E87F4C2E0279ED2E5C1C8BA886351502A1EF3859A79818D668FE7BEA919D103D84FBC8415A440DCCC88B020C4B42EA5F74401CD257D7936B62808FBF7D66725B85F465E23; 
        c2[0] = 2048'h02C12492280C084C4303DB5C6DF211274C244D704A4471ACC8049A4F0CE13A3B60AC47F58938AEE577E09EAB6B8245AB1A0F1BBC80601A51DADC547EC54327821E720617FE8F91E18A4EA008F2248763C14DD97C63935E051E91DF7D97FAA731B5459AAE150E9CBD467CAE9313359F243694D0C1CF4D4F05AE88AC5FFDFAB62EA5444C4F62D749B34C7A2FC4DC375CA7EC24A1CB2FBE19097CD46AF8D1A1BB361B36DE39C4FA14048B0A2DBD5BCA260336B57262CE024912161F43B6FB5A9C3285B531CF510F66FBC7A5FE0C88122AB1CBF7CFF1A2A5BD87534B4CDCDF7CF0D39C5CB26637F9E16D93CD261007424C24187E3C062EFB2D6BB3A687A77F3513B2;
		r2[0] = 256'hB11E4C9D9DD54B52ED1160846A0C6FF2B0E62B5DABFFD41B643188DE92A775E4;		
		//TEST VECTOR OUTPUT 0
		m[0] = 256'hDE8F939E96918B9A878B8B9A8C8BDEDEDE8F939E96918B9A878B8B9A8C8BDEDE;
		
		
		//TEST VECTOR INPUT 1
		c1[1]=2048'hABD2CD28588EDE0CD8C7E3686229C1253764BF347B1DAA1EC369F2671D3AE1FA08929B4F4B785D6AA8F5F7CF6536989719F258CE16A9129A1C03FF4DC368D50645E9DECBB75CA8057CF7DB12E21C28BD4EEE18D22A2AD124C3BB8D80C4CCCD65AB3D005DEB7FC949BEA0F0823D9E1CED76117DC2549E028589199DDC07AEAB53A2B53416389C36A42ACE51B277E288D07FABE78D45A344EF21E5D5349957C109512DD9A7C1B5F0D757A9844D0834E7CBDCCD7EC02E018E04396E809E87F4C2E0279ED2E5C1C8BA886351502A1EF3859A79818D668FE7BEA919D103D84FBC8415A440DCCC88B020C4B42EA5F74401CD257D7936B62808FBF7D66725B85F465E23; 
        c2[1] = 2048'h02C12492280C084C4303DB5C6DF211274C244D704A4471ACC8049A4F0CE13A3B60AC47F58938AEE577E09EAB6B8245AB1A0F1BBC80601A51DADC547EC54327821E720617FE8F91E18A4EA008F2248763C14DD97C63935E051E91DF7D97FAA731B5459AAE150E9CBD467CAE9313359F243694D0C1CF4D4F05AE88AC5FFDFAB62EA5444C4F62D749B34C7A2FC4DC375CA7EC24A1CB2FBE19097CD46AF8D1A1BB361B36DE39C4FA14048B0A2DBD5BCA260336B57262CE024912161F43B6FB5A9C3285B531CF510F66FBC7A5FE0C88122AB1CBF7CFF1A2A5BD87534B4CDCDF7CF0D39C5CB26637F9E16D93CD261007424C24187E3C062EFB2D6BB3A687A77F3513B2;
		r2[1] = 256'h5555555555555555555555555555555555555555555555555555555555555555;
		//TEST VECTOR OUTPUT 1
		m[1]=256'h4A1F9A9F2DD5F6E178A873CCD99C5652ECC6083544EE9FC7CC78A4C8E8B01342;

		
		//TEST_VECTOR INPUT 2
		c1[2]=2048'h9DB7F7ECAFFEB4AEA00FA4A7EE521BCAE8132BEDC84A66DE3A1E9038AC7BB97B2905727713F5F83EE8F627DF67E39AEFE8602BA617A1C8525018B1916D7B022455297EE9DFA4B7F21AEC05D22387775784A14F4B501263873C2026FA4366D16CF4038A3E65B01044A8388B2B9CF62FC9A05A0DCB2CB6D442C6F6ACBF7DBCAEB41B98DE20FC39F1D3910BA2178638EB46F05D5AE95905403D2E47786E0451C6EC8AD70F03170FCC6768393A2113BCBB8D0B66CE2062C55A1558A0F1B5C182CF3F44B68DAF28E72EE190F2801FCA1F2A728BEA639D82A68AC57DF9AB761D17A5E66AFADC5D2E0C652437EC8F6F443A4B39767E29D71F31BD9E2CC8322E3CB7C379; 
        c2[2] = 2048'h4D9AB5CF42CD447F843E6696161A8042AE71009FEDCEC6393D3E3065DA36E87F281622AA857BF7A93AAA52E0CA27871148EF80CAB7248C7FD37C92049CDEA44D56E76D00F8D6BC33795764427BE66E16B61E1DEAB61DC70389A3D609E8F30C5C050489E3B9871971334D5160C04A03ED0D7C4D7DC0BA97391F69765400B34A864A083C765C8B5C2E04ACB769CC67433F9FE8FB6CA58E9B4B6D50C45011C4717F02CA15B80D8D91821F1F7914032D6DB72636B517B7DDE1BC6CF1080BC70C1D403A376601518B311257794D861586473FE30C29DA0F5AC825E9594B1C8485BB120238DACCC76B669A04A2BF3D8F5AA6E5A9C828BAE24230E06E4118F840158ED1;
		r2[2] = 256'h5555555555555555555555555555555555555555555555555555555555555555;
		//TEST VECTOR OUTPUT 2
		m[2]=256'h8836C88E4A4F60FE209DB95E997147F9CED1D3B2EFC6980E7939FE9BB5472482;
		
		//TEST_VECTOR INPUT 3
		c1[3]=2048'hBE3A84DCAC7B7878A68FD66D9A8A958EB26573BB5D0030BF08F95D85526D5AEF14EE7F55D6CA382E50B014536CC345E3AB8A46DAA2D374BD0AC4D4B31DF3253834E658AC0B40B7E72D446BADEBDC5344B37AD9C726804D4079C14A12F685105D8ADC1E856A99D86BD25EAD5D68C7D22D708FFFA3195E12B499183249F5A5F1A7330E220FBECEDA1AA16DF4C8D3EFD8B1EF1DA166866D432CC96AEB52668F762D6C05295AA4C26FA2B5E401AB694AE1AA3F8059D8048B20C6CAF64553E387B312F7C75BCDC57E0D2CADFFB1A16C98C27F894012E6359E28E1E5638FAD7D1BBE2D31EFB4A1EE13E4C0732C2A05D97E5A3233C5CAA275CDDC589F7AE762EE5FAF92; 
        c2[3] = 2048'h4084707CE32190755C52720973230766085D79B7501CB864125B02742B81D1147D98C4550EDD4E12345545225AD3E57B72815991E5F74124CC0C6A881F1B49DA805E8BDB5FB1582B0E6782FBD695093E768602AA27402E85569F890273C5F2180B6BA2FC47091CC0282E837D74464E36022B1299199EB2402F0685BF2856B8487469EF6BF20DF76D694181F9BCB010105152FF47B359FF6DB862CC41835D98D2753A090A56E344F534A52FD81CB9837EF5756DD55670951A6A82B28F40B5E90CA9AF8382A705B96E0E0A130E2A2750FEDF4D4B0EEFC27B04A5EEA0D430B5B47EBB222E6D3500D6F0BBFFC74C5D86F04331B3AFF26ADA1CE6337FDDB965E43D58;
		r2[3] = 256'h3F1C77C5A86E5AF119A4073F51FDAEA7489DB4B3F3172961CC2BCB4ED2E28EB7;
		//TEST VECTOR OUTPUT 3
		m[3]=256'hE258A9A14BF88AF77E50CFE0A27F35EE8C041F0AB7C52FBBCDC7328F93AD56FB;
		
		
		//TEST_VECTOR INPUT 4
		c1[4]=2048'h55955207F8E3C9DF775B52F0FA2FA71EFE5CA27C05C213E1064739B6231D8AD7C16EF7C834E84B4EEAD07B0F882CEC04D7BEBB0842C15393817101B0A913BC5AD07B2F8B38DFEA1511539134460458DA5B35DE64618294FF1B6346C3E69AA5D714213E0CFC60CBF8D4A5F6EE2F1E4C7C182754733457F84EE62F70D498262E77AEBA2025C64CDDFB69E58FBB8BA6D0FC17C9AABF4532A2BC28EF26CDEFF760AD777F3F75FD27B6CC4A59094FC73DC3405F74BDCE7B6F317B1764FCD6260F0C7285E2440B665BFEEF13DE74EC2853F4EB2CE66E7B3A9231074EC45D992ADFA63A4C97CAE5F8B7D90375CDBA9DFA4453C46F11A940A19137F2B03CBDA2FD64C433; 
        c2[4] = 2048'h383A9F91890FF2750C6A056DD7940C0A70982A19366699BB5FD735BBFA360510088764C0A4C13A5F1E3433368BCA1B1B30B331653AABFDD2A0E432B2DA367BD564F4644F304C65AF5ECAFB0132623094BB198B4605A0D65D89911FC08E8885E7B95DD29766CBEAE34D81066FB0FBA03EB39EF6C0AA34D0C31D07C69E2CA521D5451348D490982EF02EA8F9839A67AC8EF1E10CF091C43D848D0E795E054BB7A860312A9CB2CBAD1B6F0691023A4C29B65A37AD4B99304380D6C346811FCFEAE2F15122693C0FDB2533F1808B323A4940E5C203CD9E6B0E2FEDA9C6EE842CFB9F1CAF11E929C0794B5C8717A8AFB84E9B7A069C5CCC1C448542F37C9349ECA107;
		r2[4] = 256'h3F1C77C5A86E5AF119A4073F51FDAEA7489DB4B3F3172961CC2BCB4ED2E28EB7;
		//TEST VECTOR OUTPUT 4
		m[4]=256'hDFF77C878F7F57D877523ACA99ADFB1FE09BE91E309D3459E575809B6106D9DF;
		
		// Initialize Inputs
		clk = 0;
		//data_rdy = 0;
		c1_in = 0;
		c2_in = 0;
		r2_in = 0;
		reset = 0;
		load = 0;
		c1_temp = 0;
		c2_temp = 0;
		r2_temp = 0;
		start=0;

		#(CLOCK_PERIOD*10);

		reset = 1;
		#(CLOCK_PERIOD);
		#(CLOCK_PERIOD);
		#(CLOCK_PERIOD);
		#(CLOCK_PERIOD);
		#(CLOCK_PERIOD);
		reset = 0;
		#(CLOCK_PERIOD);
		#(CLOCK_PERIOD);
		#(CLOCK_PERIOD);

		//main test loop
		for (j=0;j<ITERATION_SIZE;j=j+1)
		begin
			
			for (i=0;i<256;i=i+1)
			begin
				//#(CLOCK_PERIOD/2);
				load = 1;
				c1_temp=c1[j]>>i*8;
				c2_temp=c2[j]>>i*8;
				r2_temp=r2[j]>>i;
				c1_in = c1_temp[7:0];
				c2_in = c2_temp[7:0];
				r2_in = r2_temp[0];
				#(CLOCK_PERIOD);
			end
			load = 0;
			#(CLOCK_PERIOD*3);
			start=1;
			#(CLOCK_PERIOD*2);
			start=0;
			
			//define a wait period here -- this depends on the execution time of your design
			// for example #(CLOCK_PERIOD*10) ;
			// your design is likely to execute more than this
          
          	// wait(dut.mult_done);
          	// $display("c1*r2: %h", dut.mem_state);
          
          	// wait(dut.add_done);
          	// $display("c1*r2 + c2: %h", dut.mem_state);
          
			// wait(dut.out_done);
          	#(CLOCK_PERIOD*99201.5);

          	// $display("time: %0t", $time);
          	// $display("message_fifo: %h", message_fifo);
          	// $display("cnt_out: %d", cnt_out);
          	// $display("cmp: %0d\n", cmp);

          	#(CLOCK_PERIOD*1.5);
		end

		$stop;
	end
	
	//generate clock
	always #(CLOCK_PERIOD/2) clk = ~clk;
    
	
	//check if output matches the expected one
	reg [255:0]message_fifo;
	reg [8:0]cnt_out;
	reg valid_d1;
	always @ (posedge clk or posedge reset)
	begin
		if (reset)
		begin
			cnt_out<=0;
			message_fifo <=0;
		end
		else if (valid)
		begin
			cnt_out<=cnt_out+1;
			message_fifo[cnt_out] <= message_out;
		end
		else if (cnt_out==256)
			cnt_out<=0;
	end
	
	//cmp should be high for one clock cycle per evaluation (right after the output is generated)
	assign cmp=(cnt_out==256 && (message_fifo == m[j]))?1:0;
  
  	// initial begin
    //   $dumpfile("dump.vcd");
    //   $dumpvars(0, dut);
    // end
endmodule
